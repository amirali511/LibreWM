module main

import librewm

pub fn main () {
	panic ("Shit! I forgot to write this file! Not for production and public use yet! Now go and have your cup of coffee!");	
}
