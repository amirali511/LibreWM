module main

import librewm

pub fn main () {
		
}
